Counter
  
